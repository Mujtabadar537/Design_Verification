interface dut_if();

logic [15:0]in1;
logic [15:0]in2;
logic cin;

logic [15:0]sum;
logic carry;


endinterface

interface dut_if();

bit clk,reset,d;
bit q,qbar;

endinterface

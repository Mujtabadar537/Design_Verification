interface dut_if();

logic in1,in2,cin;
logic sum,cout;


endinterface

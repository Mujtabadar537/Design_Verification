interface design_interface(input logic clk , reset);

logic in;
logic out;

endinterface
